{"location_units": ["deg", "deg"], "location": [-117.0, 34.0]}