{"location_units": ["deg", "deg"], "location": [-112.0, 34.0]}